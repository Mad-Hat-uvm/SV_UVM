interface not_if();
    logic in;
    logic out;
endinterface