class scoreboard extends uvm_scoreboard;
    `uvm_component_utils(scoreboard)

    uvm_analysis_imp #(seq_item, scoreboard) item_collect_export;

    function new(string name="env", uvm_component parent=null);
        super.new(name, parent);

        item_collect_export = new("item_collect_export", this);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
    endfunction

    function void write(seq_item req);
        $display("--------------------------------------------------------");

        if(req.out == ~req.in) begin
        `uvm_info(get_type_name(), $sformatf("MATCH IN=%0d, OUT=%0d", req.in, req.out), UVM_LOW);
        end

        else begin
            `uvm_info(get_type_name(), $sformatf("NOT MATCH IN=%0d, OUT=%0d", req.in, req.out), UVM_LOW);  
        end

        $display("--------------------------------------------------------");
    endfunction
endclass