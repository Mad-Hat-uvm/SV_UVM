interface add_if(
  input logic clk,
  input logic reset
);

  logic [7:0] ip1;
  logic [7:0] ip2;
  logic [8:0] out;
  
endinterface
