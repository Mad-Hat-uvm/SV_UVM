`include "transaction.sv"

`include "read_data.sv"

`include "read_err.sv"

`include "reset_dut.sv"

`include "write_data.sv"

`include "write_err.sv"

`include "write_read.sv"

`include "writeb_readb.sv"

`include "driver.sv"

`include "mon.sv"

`include "sco.sv"

`include "agent.sv"

`include "env.sv"

`include "apb_config.sv"

`include "test.sv"