`include "seq_item.sv"

`include "base_seq.sv"

`include "driver.sv"

`include "monitor.sv"

`include "scoreboard.sv"

`include "active_agent.sv"

`include "env.sv"
